// SPDX-FileCopyrightText: 2024 Ayuub Mohamud <ayuub.mohamud@outlook.com>
// SPDX-License-Identifier: CERN-OHL-W-2.0

//  -----------------------------------------------------------------------------------------
//  | Copyright (C) Ayuub Mohamud 2024.                                                     |
//  |                                                                                       |
//  | This source describes Open Hardware (RTL) and is licensed under the CERN-OHL-W v2.    |
//  |                                                                                       |
//  | You may redistribute and modify this source and make products using it under          |
//  | the terms of the CERN-OHL-W v2 (https://ohwr.org/cern_ohl_w_v2.txt).                  |
//  |                                                                                       |
//  | This source is distributed WITHOUT ANY EXPRESS OR IMPLIED WARRANTY,                   |
//  | INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY AND FITNESS FOR A                  |
//  | PARTICULAR PURPOSE. Please see the CERN-OHL-W v2 for applicable conditions.           |
//  |                                                                                       |
//  | Source location: https://github.com/AyuubMohamud/Biriq                                |
//  |                                                                                       |
//  | As per CERN-OHL-W v2 section 4, should You produce hardware based on this             |
//  | source, You must where practicable maintain the Source Location visible               |
//  | in the same manner as is done within this source.                                     |
//  |                                                                                       |
//  -----------------------------------------------------------------------------------------
module engine (
    input  wire         core_clock_i,
    output wire         dcache_flush_o,
    input  wire         dcache_flush_resp,
    input  wire         ins0_port_i,
    input  wire         ins0_dnagn_i,
    input  wire  [ 6:0] ins0_alu_type_i,
    input  wire  [ 6:0] ins0_alu_opcode_i,
    input  wire         ins0_alu_imm_i,
    input  wire  [ 5:0] ins0_ios_type_i,
    input  wire  [ 2:0] ins0_ios_opcode_i,
    input  wire  [ 3:0] ins0_special_i,
    input  wire  [ 4:0] ins0_rs1_i,
    input  wire  [ 4:0] ins0_rs2_i,
    input  wire  [ 4:0] ins0_dest_i,
    input  wire  [31:0] ins0_imm_i,
    input  wire  [ 2:0] ins0_reg_props_i,
    input  wire         ins0_dnr_i,
    input  wire         ins0_mov_elim_i,
    input  wire  [ 1:0] ins0_hint_i,
    input  wire         ins0_excp_valid_i,
    input  wire  [ 3:0] ins0_excp_code_i,
    input  wire         ins1_port_i,
    input  wire         ins1_dnagn_i,
    input  wire  [ 6:0] ins1_alu_type_i,
    input  wire  [ 6:0] ins1_alu_opcode_i,
    input  wire         ins1_alu_imm_i,
    input  wire  [ 5:0] ins1_ios_type_i,
    input  wire  [ 2:0] ins1_ios_opcode_i,
    input  wire  [ 3:0] ins1_special_i,
    input  wire  [ 4:0] ins1_rs1_i,
    input  wire  [ 4:0] ins1_rs2_i,
    input  wire  [ 4:0] ins1_dest_i,
    input  wire  [31:0] ins1_imm_i,
    input  wire  [ 2:0] ins1_reg_props_i,
    input  wire         ins1_dnr_i,
    input  wire         ins1_mov_elim_i,
    input  wire  [ 1:0] ins1_hint_i,
    input  wire         ins1_excp_valid_i,
    input  wire  [ 3:0] ins1_excp_code_i,
    input  wire         ins1_valid_i,
    input  wire  [29:0] insbundle_pc_i,
    input  wire  [ 1:0] btb_btype_i,
    input  wire  [ 1:0] btb_bm_pred_i,
    input  wire  [29:0] btb_target_i,
    input  wire         btb_vld_i,
    input  wire         btb_idx_i,
    input  wire         btb_way_i,
    input  wire         valid_i,
    output wire         rn_busy_o,
    output wire  [ 6:0] ms_ins0_opcode_o,
    output wire  [ 6:0] ms_ins0_ins_type,
    output wire         ms_ins0_imm_o,
    output wire  [31:0] ms_ins0_immediate_o,
    output wire  [ 5:0] ms_ins0_dest_o,
    output wire  [ 1:0] ms_ins0_hint_o,
    output wire         ms_ins0_valid,
    output wire  [ 6:0] ms_ins1_opcode_o,
    output wire  [ 6:0] ms_ins1_ins_type,
    output wire         ms_ins1_imm_o,
    output wire  [31:0] ms_ins1_immediate_o,
    output wire  [ 5:0] ms_ins1_dest_o,
    output wire  [ 1:0] ms_ins1_hint_o,
    output wire         ms_ins1_valid,
    output wire  [ 3:0] ms_pack_id,
    output wire  [29:0] ms_rn_pc_o,
    output wire  [ 1:0] ms_rn_bm_pred_o,
    output wire  [ 1:0] ms_rn_btype_o,
    output wire         ms_rn_btb_vld_o,
    output wire  [29:0] ms_rn_btb_target_o,
    output wire         ms_rn_btb_way_o,
    output wire         ms_rn_btb_idx_o,
    output wire  [ 3:0] ms_rn_btb_pack,
    output wire         ms_rn_btb_wen,
    output wire  [17:0] ms_p0_data_o,
    output wire         ms_p0_sc_o,
    output wire         ms_p0_mc_o,
    output wire         ms_p0_vld_o,
    output wire         ms_p0_rs1_vld_o,
    output wire         ms_p0_rs2_vld_o,
    output wire         ms_p0_rs1_rdy,
    output wire         ms_p0_rs2_rdy,
    output wire  [17:0] ms_p1_data_o,
    output wire         ms_p1_sc_o,
    output wire         ms_p1_mc_o,
    output wire         ms_p1_vld_o,
    output wire         ms_p1_rs1_vld_o,
    output wire         ms_p1_rs2_vld_o,
    output wire         ms_p1_rs1_rdy,
    output wire         ms_p1_rs2_rdy,
    input  wire         ms_p0_busy_i,
    input  wire         ms_p1_busy_i,
    // memory Sys  
    output wire         memSys_renamer_pkt_vld_o,
    output wire  [ 5:0] memSys_pkt0_rs1_o,
    output wire  [ 5:0] memSys_pkt0_rs2_o,
    output wire  [ 5:0] memSys_pkt0_dest_i,
    output wire  [31:0] memSys_pkt0_immediate_o,
    output wire  [ 5:0] memSys_pkt0_ios_type_o,
    output wire  [ 2:0] memSys_pkt0_ios_opcode_o,
    output wire  [ 4:0] memSys_pkt0_rob_o,
    output wire         memSys_pkt0_vld_o,
    output wire  [ 5:0] memSys_pkt1_rs1_o,
    output wire  [ 5:0] memSys_pkt1_rs2_o,
    output wire  [ 5:0] memSys_pkt1_dest_o,
    output wire  [31:0] memSys_pkt1_immediate_o,
    output wire  [ 5:0] memSys_pkt1_ios_type_o,
    output wire  [ 2:0] memSys_pkt1_ios_opcode_o,
    output wire         memSys_pkt1_vld_o,
    input  wire         memSys_full,
    input  wire         cpm,
    input  wire         mie,
    input  wire  [ 2:0] machine_interrupts,
    input  wire  [ 4:0] alu0_rob_slot_i,
    input  wire         alu0_rob_complete_i,
    input  wire         alu0_call_i,
    input  wire         alu0_ret_i,
    input  wire  [ 4:0] alu1_rob_slot_i,
    input  wire         alu1_rob_complete_i,
    input  wire  [ 4:0] agu0_rob_slot_i,
    input  wire         agu0_rob_complete_i,
    input  wire  [ 4:0] ldq_rob_slot_i,
    input  wire         ldq_rob_complete_i,
    input  wire         alu0_reg_ready,
    input  wire  [ 5:0] alu0_reg_dest,
    input  wire         alu1_reg_ready,
    input  wire  [ 5:0] alu1_reg_dest,
    input  wire         alul_reg_ready,
    input  wire  [ 5:0] alul_reg_dest,
    output wire         stb_c0,
    output wire         stb_c1,
    input  wire         stb_emp,
    input  wire         alu_excp_i,
    input  wire  [ 4:0] alu_excp_code_i,
    input  wire  [ 5:0] rob_i,
    input  wire  [29:0] c1_btb_vpc_i,
    input  wire  [29:0] c1_btb_target_i,
    input  wire  [ 1:0] c1_cntr_pred_i,
    input  wire         c1_bnch_tkn_i,
    input  wire  [ 1:0] c1_bnch_type_i,
    input  wire         c1_bnch_present_i,
    input  wire  [ 5:0] completed_rob_id,
    input  wire  [ 4:0] exception_code_i,
    input  wire  [31:0] exception_addr,
    input  wire         exception_i,
    input  wire         icache_idle,
    input  wire         mem_block_i,
    output wire         icache_flush,
    output wire         flush,
    output       [29:0] flush_address,
    output wire         rcu_block,
    output wire  [ 4:0] oldest_instruction,
    output wire         rename_flush_o,
    output wire         ins_commit0,
    output wire         ins_commit1,
    output wire         mret,
    output wire         take_exception,
    output wire         take_interrupt,
    output wire  [29:0] tmu_epc_o,
    output wire  [31:0] tmu_mtval_o,
    output wire  [ 3:0] tmu_mcause_o,
    input  wire  [29:0] mepc_i,
    input  wire  [31:0] mtvec_i,
    output wire  [29:0] c1_btb_vpc_o,
    output wire  [29:0] c1_btb_target_o,
    output wire  [ 1:0] c1_cntr_pred_o,
    output wire         c1_bnch_tkn_o,
    output wire  [ 1:0] c1_bnch_type_o,
    output wire         c1_btb_mod_o,
    output wire         c1_call_affirm_o,
    output wire         c1_ret_affirm_o,
    input  wire         p0_we_i,
    input  wire  [31:0] p0_we_data,
    input  wire  [ 5:0] p0_we_dest,
    input  wire         p0_ex_i,
    input  wire  [31:0] p0_ex_data,
    input  wire  [ 5:0] p0_ex_dest,
    input  wire         p1_we_i,
    input  wire  [31:0] p1_we_data,
    input  wire  [ 5:0] p1_we_dest,
    input  wire         p1_ex_i,
    input  wire  [31:0] p1_ex_data,
    input  wire  [ 5:0] p1_ex_dest,
    input  wire         p2_we_i,
    input  wire  [31:0] p2_we_data,
    input  wire  [ 5:0] p2_we_dest,
    input  wire  [ 5:0] p0_rd_src,
    output logic [31:0] p0_rd_datas,
    input  wire  [ 5:0] p1_rd_src,
    output logic [31:0] p1_rd_datas,
    input  wire  [ 5:0] p2_rd_src,
    output logic [31:0] p2_rd_datas,
    input  wire  [ 5:0] p3_rd_src,
    output logic [31:0] p3_rd_datas,
    input  wire  [ 5:0] p4_rd_src,
    output logic [31:0] p4_rd_datas,
    input  wire  [ 5:0] p5_rd_src,
    output logic [31:0] p5_rd_datas,
    input  wire  [ 5:0] r4_vec_indx,
    output wire         r4,
    input  wire  [ 5:0] r5_vec_indx,
    output wire         r5
);
  wire rename_flush = flush;
  reg [5:0] c0 = 6'd0;
  reg [5:0] c1 = 6'd1;
  reg [5:0] c2 = 6'd2;
  reg [5:0] c3 = 6'd3;
  always_ff @(posedge core_clock_i) begin
    if (rename_flush) begin
      c0 <= c0 + 4;
      c1 <= c1 + 4;
      c2 <= c2 + 4;
      c3 <= c3 + 4;
    end
  end
  irf integerRegisterFile (
      core_clock_i,
      p0_we_i,
      p0_we_data,
      p0_we_dest,
      p0_ex_i,
      p0_ex_data,
      p0_ex_dest,
      p1_we_i,
      p1_we_data,
      p1_we_dest,
      p1_ex_i,
      p1_ex_data,
      p1_ex_dest,
      p2_we_i,
      p2_we_data,
      p2_we_dest,
      p0_rd_src,
      p0_rd_datas,
      p1_rd_src,
      p1_rd_datas,
      p2_rd_src,
      p2_rd_datas,
      p3_rd_src,
      p3_rd_datas,
      p4_rd_src,
      p4_rd_datas,
      p5_rd_src,
      p5_rd_datas
  );
  wire [5:0] p0_vec_indx;
  wire       p0_busy_vld;
  wire [5:0] p1_vec_indx;
  wire       p1_free_vld = 1'b0;
  wire       p1_busy_vld;
  wire [5:0] p2_vec_indx = rename_flush ? c0 : alu0_reg_dest;
  wire       p2_free_vld = rename_flush | alu0_reg_ready;  // early wake
  wire [5:0] p3_vec_indx = rename_flush ? c1 : alu1_reg_dest;
  wire       p3_free_vld = rename_flush | alu1_reg_ready;
  wire [5:0] p4_vec_indx = rename_flush ? c2 : p2_we_dest;
  wire       p4_free_vld = rename_flush | p2_we_i;
  wire [5:0] p5_vec_indx = rename_flush ? c3 : alul_reg_dest;
  wire       p5_free_vld = rename_flush | alul_reg_ready;
  wire [5:0] r0_vec_indx;
  wire       r0;
  wire [5:0] r1_vec_indx;
  wire       r1;
  wire [5:0] r2_vec_indx;
  wire       r2;
  wire [5:0] r3_vec_indx;
  wire       r3;
  rst rst (
      core_clock_i,
      p0_vec_indx,
      p0_busy_vld,
      p1_vec_indx,
      p1_free_vld,
      p1_busy_vld,
      p2_vec_indx,
      p2_free_vld,
      p3_vec_indx,
      p3_free_vld,
      p4_vec_indx,
      p4_free_vld,
      p5_vec_indx,
      p5_free_vld,
      r0_vec_indx,
      r0,
      r1_vec_indx,
      r1,
      r2_vec_indx,
      r2,
      r3_vec_indx,
      r3,
      r4_vec_indx,
      r4,
      r5_vec_indx,
      r5
  );
  wire        i_wr_en0;
  wire  [5:0] i_wr_data0;
  wire        o_full0;
  wire        i_wr_en1;
  wire  [5:0] i_wr_data1;
  wire        o_full1;
  wire        i_rd0;
  logic [5:0] o_rd_data0;
  wire        o_empty0;
  wire        i_rd1;
  logic [5:0] o_rd_data1;
  wire        o_empty1;
  freelist freelist (
      core_clock_i,
      i_wr_en0,
      i_wr_data0,
      o_full0,
      i_wr_en1,
      i_wr_data1,
      o_full1,
      i_rd0,
      o_rd_data0,
      o_empty0,
      i_rd1,
      o_rd_data1,
      o_empty1
  );
  wire [4:0] rob0_status;
  wire       commit0;
  wire       rob0_status_o;
  wire       rob0_call_o;
  wire       rob0_ret_o;
  wire [4:0] rob1_status;
  wire       commit1;
  wire       rob1_status_o;
  wire       rob1_call_o;
  wire       rob1_ret_o;
  ciff ciff (
      core_clock_i,
      flush,
      alu0_rob_slot_i,
      alu0_rob_complete_i,
      alu0_call_i,
      alu0_ret_i,
      alu1_rob_slot_i,
      alu1_rob_complete_i,
      agu0_rob_slot_i,
      agu0_rob_complete_i,
      ldq_rob_slot_i,
      ldq_rob_complete_i,
      rob0_status,
      commit0,
      rob0_status_o,
      rob0_call_o,
      rob0_ret_o,
      rob1_status,
      commit1,
      rob1_status_o,
      rob1_call_o,
      rob1_ret_o
  );
  wire [29:0] packet_pc;
  wire        ins0_is_mov_elim;
  wire        ins0_register_allocated;
  wire [ 4:0] ins0_arch_reg;
  wire [ 5:0] ins0_old_preg;
  wire [ 5:0] ins0_new_preg;
  wire [ 3:0] ins0_excp_code;
  wire        ins0_excp_valid;
  wire [ 3:0] ins0_special;
  wire        ins0_is_store;
  wire        ins1_is_mov_elim;
  wire        ins1_register_allocated;
  wire [ 4:0] ins1_arch_reg;
  wire [ 5:0] ins1_old_preg;
  wire [ 5:0] ins1_new_preg;
  wire [ 3:0] ins1_excp_code;
  wire        ins1_excp_valid;
  wire [ 3:0] ins1_special;
  wire        ins1_is_store;
  wire        ins1_valid;
  wire        push_packet;
  wire        rcu_busy;
  wire [ 4:0] rcu_pack;
  wire [ 4:0] arch_reg0;
  wire [ 4:0] arch_reg1;
  wire [ 5:0] phys_reg0;
  wire [ 5:0] phys_reg1;

  rename renamer (
      core_clock_i,
      rename_flush_o,
      flush,
      ins0_port_i,
      ins0_dnagn_i,
      ins0_alu_type_i,
      ins0_alu_opcode_i,
      ins0_alu_imm_i,
      ins0_ios_type_i,
      ins0_ios_opcode_i,
      ins0_special_i,
      ins0_rs1_i,
      ins0_rs2_i,
      ins0_dest_i,
      ins0_imm_i,
      ins0_reg_props_i,
      ins0_dnr_i,
      ins0_mov_elim_i,
      ins0_hint_i,
      ins0_excp_valid_i,
      ins0_excp_code_i,
      ins1_port_i,
      ins1_dnagn_i,
      ins1_alu_type_i,
      ins1_alu_opcode_i,
      ins1_alu_imm_i,
      ins1_ios_type_i,
      ins1_ios_opcode_i,
      ins1_special_i,
      ins1_rs1_i,
      ins1_rs2_i,
      ins1_dest_i,
      ins1_imm_i,
      ins1_reg_props_i,
      ins1_dnr_i,
      ins1_mov_elim_i,
      ins1_hint_i,
      ins1_excp_valid_i,
      ins1_excp_code_i,
      ins1_valid_i,
      insbundle_pc_i,
      btb_btype_i,
      btb_bm_pred_i,
      btb_target_i,
      btb_vld_i,
      btb_idx_i,
      btb_way_i,
      valid_i,
      rn_busy_o,
      packet_pc,
      ins0_is_mov_elim,
      ins0_register_allocated,
      ins0_arch_reg,
      ins0_old_preg,
      ins0_new_preg,
      ins0_excp_code,
      ins0_excp_valid,
      ins0_special,
      ins0_is_store,
      ins1_is_mov_elim,
      ins1_register_allocated,
      ins1_arch_reg,
      ins1_old_preg,
      ins1_new_preg,
      ins1_excp_code,
      ins1_excp_valid,
      ins1_special,
      ins1_is_store,
      ins1_valid,
      push_packet,
      rcu_busy,
      rcu_pack,
      arch_reg0,
      arch_reg1,
      phys_reg0,
      phys_reg1,
      ms_ins0_opcode_o,
      ms_ins0_ins_type,
      ms_ins0_imm_o,
      ms_ins0_immediate_o,
      ms_ins0_dest_o,
      ms_ins0_hint_o,
      ms_ins0_valid,
      ms_ins1_opcode_o,
      ms_ins1_ins_type,
      ms_ins1_imm_o,
      ms_ins1_immediate_o,
      ms_ins1_dest_o,
      ms_ins1_hint_o,
      ms_ins1_valid,
      ms_pack_id,
      ms_rn_pc_o,
      ms_rn_bm_pred_o,
      ms_rn_btype_o,
      ms_rn_btb_vld_o,
      ms_rn_btb_target_o,
      ms_rn_btb_way_o,
      ms_rn_btb_idx_o,
      ms_rn_btb_pack,
      ms_rn_btb_wen,
      ms_p0_data_o,
      ms_p0_sc_o,
      ms_p0_mc_o,
      ms_p0_vld_o,
      ms_p0_rs1_vld_o,
      ms_p0_rs2_vld_o,
      ms_p0_rs1_rdy,
      ms_p0_rs2_rdy,
      ms_p1_data_o,
      ms_p1_sc_o,
      ms_p1_mc_o,
      ms_p1_vld_o,
      ms_p1_rs1_vld_o,
      ms_p1_rs2_vld_o,
      ms_p1_rs1_rdy,
      ms_p1_rs2_rdy,
      ms_p0_busy_i,
      ms_p1_busy_i,
      memSys_renamer_pkt_vld_o,
      memSys_pkt0_rs1_o,
      memSys_pkt0_rs2_o,
      memSys_pkt0_dest_i,
      memSys_pkt0_immediate_o,
      memSys_pkt0_ios_type_o,
      memSys_pkt0_ios_opcode_o,
      memSys_pkt0_rob_o,
      memSys_pkt0_vld_o,
      memSys_pkt1_rs1_o,
      memSys_pkt1_rs2_o,
      memSys_pkt1_dest_o,
      memSys_pkt1_immediate_o,
      memSys_pkt1_ios_type_o,
      memSys_pkt1_ios_opcode_o,
      memSys_pkt1_vld_o,
      memSys_full,
      p0_vec_indx,
      p0_busy_vld,
      p1_vec_indx,
      p1_busy_vld,
      r0_vec_indx,
      r0,
      r1_vec_indx,
      r1,
      r2_vec_indx,
      r2,
      r3_vec_indx,
      r3,
      i_rd0,
      o_rd_data0,
      o_empty0,
      i_rd1,
      o_rd_data1,
      o_empty1
  );
  retireControlUnit rcu0 (
      core_clock_i,
      dcache_flush_o,
      dcache_flush_resp,
      cpm,
      mie,
      machine_interrupts,
      packet_pc,
      ins0_is_mov_elim,
      ins0_register_allocated,
      ins0_arch_reg,
      ins0_old_preg,
      ins0_new_preg,
      ins0_excp_code,
      ins0_excp_valid,
      ins0_special,
      ins0_is_store,
      ins1_is_mov_elim,
      ins1_register_allocated,
      ins1_arch_reg,
      ins1_old_preg,
      ins1_new_preg,
      ins1_excp_code,
      ins1_excp_valid,
      ins1_special,
      ins1_is_store,
      ins1_valid,
      push_packet,
      rcu_busy,
      rcu_pack,
      arch_reg0,
      arch_reg1,
      phys_reg0,
      phys_reg1,
      rob0_status,
      commit0,
      rob0_status_o,
      rob0_call_o,
      rob0_ret_o,
      rob1_status,
      commit1,
      rob1_status_o,
      rob1_call_o,
      rob1_ret_o,
      stb_c0,
      stb_c1,
      stb_emp,
      i_wr_en0,
      i_wr_data0,
      i_wr_en1,
      i_wr_data1,
      alu_excp_i,
      alu_excp_code_i,
      rob_i,
      c1_btb_vpc_i,
      c1_btb_target_i,
      c1_cntr_pred_i,
      c1_bnch_tkn_i,
      c1_bnch_type_i,
      c1_bnch_present_i,
      completed_rob_id,
      exception_code_i,
      exception_addr,
      exception_i,
      icache_idle,
      mem_block_i,
      icache_flush,
      flush,
      flush_address,
      rcu_block,
      oldest_instruction,
      rename_flush_o,
      ins_commit0,
      ins_commit1,
      mret,
      take_exception,
      take_interrupt,
      tmu_epc_o,
      tmu_mtval_o,
      tmu_mcause_o,
      mepc_i,
      mtvec_i,
      c1_btb_vpc_o,
      c1_btb_target_o,
      c1_cntr_pred_o,
      c1_bnch_tkn_o,
      c1_bnch_type_o,
      c1_btb_mod_o,
      c1_call_affirm_o,
      c1_ret_affirm_o
  );
endmodule
