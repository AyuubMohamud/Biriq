module ixu (

  );

endmodule
