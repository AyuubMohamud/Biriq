localparam UIB_JAL = 3'd0;
localparam UIB_JALR = 3'd1;
localparam UIB_AUIPC = 3'd2;
localparam UIB_OP = 3'd3;
localparam UIB_BRANCH = 3'd4;
localparam UIB_MEMORY = 3'd5;
localparam UIB_MULDIV = 3'd6;
localparam UIB_CSR = 3'd7;
localparam MEMOP_LOAD = 3'd0;
localparam MEMOP_LR = 3'd1;
localparam MEMOP_STORE = 3'd2;
localparam MEMOP_SC = 3'd3;
localparam MEMOP_AMO = 3'd4;
localparam MEMOP_CMO = 3'd5;
localparam MEMSZ_BYTE = 2'd0;
localparam MEMSZ_HALF = 2'd1;
localparam MEMSZ_WORD = 2'd2;
