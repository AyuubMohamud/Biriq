module ieu (
    
);
    
endmodule
