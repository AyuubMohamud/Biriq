// SPDX-FileCopyrightText: 2024 Ayuub Mohamud <ayuub.mohamud@outlook.com>
// SPDX-License-Identifier: CERN-OHL-W-2.0

//  -----------------------------------------------------------------------------------------
//  | Copyright (C) Ayuub Mohamud 2024.                                                     |
//  |                                                                                       |
//  | This source describes Open Hardware (RTL) and is licensed under the CERN-OHL-W v2.    |
//  |                                                                                       |
//  | You may redistribute and modify this source and make products using it under          |
//  | the terms of the CERN-OHL-W v2 (https://ohwr.org/cern_ohl_w_v2.txt).                  |
//  |                                                                                       |
//  | This source is distributed WITHOUT ANY EXPRESS OR IMPLIED WARRANTY,                   |
//  | INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY AND FITNESS FOR A                  |
//  | PARTICULAR PURPOSE. Please see the CERN-OHL-W v2 for applicable conditions.           |
//  |                                                                                       |
//  | Source location: https://github.com/AyuubMohamud/Biriq                                |
//  |                                                                                       |
//  | As per CERN-OHL-W v2 section 4, should You produce hardware based on this             |
//  | source, You must where practicable maintain the Source Location visible               |
//  | in the same manner as is done within this source.                                     |
//  |                                                                                       |
//  -----------------------------------------------------------------------------------------
// RCU
/**
**/
module retireControlUnit (
    input  wire logic cpu_clock_i,
    output wire logic dcache_flush_o,
    input  wire logic dcache_flush_resp,

    input wire logic       cpm,
    input wire logic       mie,
    input wire logic [2:0] machine_interrupts,

    input  wire logic [29:0] packet_pc,
    input  wire logic        ins0_is_mov_elim,
    input  wire logic        ins0_register_allocated,
    input  wire logic [ 4:0] ins0_arch_reg,
    input  wire logic [ 5:0] ins0_old_preg,
    input  wire logic [ 5:0] ins0_new_preg,
    input  wire logic [ 3:0] ins0_excp_code,
    input  wire logic        ins0_excp_valid,
    input  wire logic [ 3:0] ins0_special,
    input  wire logic        ins0_is_store,
    input  wire logic        ins1_is_mov_elim,
    input  wire logic        ins1_register_allocated,
    input  wire logic [ 4:0] ins1_arch_reg,
    input  wire logic [ 5:0] ins1_old_preg,
    input  wire logic [ 5:0] ins1_new_preg,
    input  wire logic [ 3:0] ins1_excp_code,
    input  wire logic        ins1_excp_valid,
    input  wire logic [ 3:0] ins1_special,
    input  wire logic        ins1_is_store,
    input  wire logic        ins1_valid,
    input  wire logic        push_packet,
    output wire logic        rcu_busy,
    output wire logic [ 4:0] rcu_pack,
    // Inst0
    input  wire logic [ 4:0] p0_logical_reg_i,
    output wire logic [ 5:0] p0_phys_reg_o,
    input  wire logic [ 4:0] p1_logical_reg_i,
    output wire logic [ 5:0] p1_phys_reg_o,
    // Inst1
    input  wire logic [ 4:0] p2_logical_reg_i,
    output wire logic [ 5:0] p2_phys_reg_o,
    input  wire logic [ 4:0] p3_logical_reg_i,
    output wire logic [ 5:0] p3_phys_reg_o,
    input  wire logic [ 4:0] p4_logical_reg_i,
    output wire logic [ 5:0] p4_phys_reg_o,
    input  wire logic [ 4:0] p5_logical_reg_i,
    output wire logic [ 5:0] p5_phys_reg_o,
    // Complete instruction bitvector
    output wire logic [ 4:0] rob0_status,
    output wire logic        commit0,
    input  wire logic        rob0_status_i,
    input  wire logic        rob0_call_i,
    input  wire logic        rob0_ret_i,
    output wire logic [ 4:0] rob1_status,
    output wire logic        commit1,
    input  wire logic        rob1_status_i,
    input  wire logic        rob1_call_i,
    input  wire logic        rob1_ret_i,
    // Store Queue/Buffer
    output wire logic        sqb_commit0,
    output wire logic        sqb_commit1,
    input  wire logic        sqb_empty,
    // free list
    output wire logic        wr_en0,
    output wire logic [ 5:0] wr_data0,
    output wire logic        wr_en1,
    output wire logic [ 5:0] wr_data1,

    // exceptions
    input wire logic        alu_excp_i,
    input wire logic [ 4:0] alu_excp_code_i,
    input wire logic [ 5:0] rob_i,
    input wire logic [29:0] c1_btb_vpc_i,
    input wire logic [29:0] c1_btb_target_i,
    input wire logic [ 1:0] c1_cntr_pred_i,
    input wire logic        c1_bnch_tkn_i,
    input wire logic [ 1:0] c1_bnch_type_i,
    input wire logic        c1_bnch_present_i,

    input wire logic [ 5:0] completed_rob_id,
    input wire logic [ 4:0] exception_code_i,
    input wire logic [31:0] exception_addr,
    input wire logic        exception_i,

    input  wire logic icache_idle,
    input  wire logic mem_block_i,
    output wire logic icache_flush,

    output wire logic        flush_o,
    output logic      [29:0] flush_address,

    output wire logic rcu_block,

    output wire logic [4:0] oldest_instruction,
    output wire logic       rename_flush_o,

    output wire logic        ins_commit0,
    output wire logic        ins_commit1,
    // exception returns
    output wire logic        mret,
    // exception handling           
    output wire logic        take_exception,
    output wire logic        take_interrupt,
    output wire logic [29:0] tmu_epc_o,
    output wire logic [31:0] tmu_mtval_o,
    output wire logic [ 3:0] tmu_mcause_o,
    input  wire logic [29:0] mepc_i,
    input  wire logic [31:0] mtvec_i,

    output wire logic [29:0] c1_btb_vpc_o,     //! SIP PC
    output wire logic [29:0] c1_btb_target_o,  //! SIP Target **if** taken
    output wire logic [ 1:0] c1_cntr_pred_o,   //! Bimodal counter prediction,
    output wire logic        c1_bnch_tkn_o,    //! Branch taken this cycle
    output wire logic [ 1:0] c1_bnch_type_o,
    output wire logic        c1_btb_mod_o,

    output wire logic c1_call_affirm_o,
    output wire logic c1_ret_affirm_o
);
  wire        full;
  wire        empty;
  wire        packet_pop;
  wire [ 4:0] rd_ptr;
  wire [ 4:0] wr_ptr;
  /*verilator lint_off UNUSEDSIGNAL*/
  wire [29:0] cpacket_pc;
  /*verilator lint_on UNUSEDSIGNAL*/
  wire        cins0_register_allocated;
  wire [ 4:0] cins0_arch_reg;
  wire [ 5:0] cins0_old_preg;
  wire [ 5:0] cins0_new_preg;
  wire [ 3:0] cins0_excp_code;
  wire        cins0_excp_valid;
  wire [ 3:0] cins0_special;
  wire        cins0_is_store;
  wire        cins1_register_allocated;
  wire [ 4:0] cins1_arch_reg;
  wire [ 5:0] cins1_old_preg;
  wire [ 5:0] cins1_new_preg;
  wire [ 3:0] cins1_excp_code;
  wire        cins1_excp_valid;
  wire [ 3:0] cins1_special;
  wire        cins1_is_store;
  wire        cins1_valid;
  wire        commit_ins0;
  wire        commit_ins1;
  wire altcommit, altcommit0, altcommit1;
  assign commit0 = commit_ins0;
  assign commit1 = commit_ins1;
  reg        partial_retire;
  reg [ 4:0] recoveryCounter0 = 5'b00000;
  reg [ 4:0] recoveryCounter1 = 5'b00001;
  reg [31:0] relavant_address;
  reg [ 4:0] exception_code;
  reg [ 5:0] exception_rob;
  reg        exception_valid = 0;
  reg [29:0] c1_btb_vpc;
  reg [29:0] c1_btb_target;
  reg [ 1:0] c1_cntr_pred;
  reg        c1_bnch_tkn;
  reg [ 1:0] c1_bnch_type;
  reg        c1_bnch_present = 0;
  localparam Normal = 3'b000;
  localparam ReclaimAndRecover = 3'b111;  // flush held high for 16 cycles
  localparam WipeInstructionCache = 3'b001;
  localparam WaitForInterrupt = 3'b010;
  localparam Await = 3'b110;
  localparam TakeInterrupt = 3'b011;
  localparam WipeDataCache = 3'b100;
  reg [2:0] retire_control_state = Normal;

  sfifospecial #(
      .DW(87)
  ) instruction_information_buffer (
      cpu_clock_i,
      1'b0,
      push_packet & !full,
      {
        packet_pc,
        ins0_register_allocated,
        ins0_arch_reg,
        ins0_old_preg,
        ins0_new_preg,
        ins0_excp_code,
        ins0_excp_valid,
        ins0_special,
        ins0_is_store,
        ins1_register_allocated,
        ins1_arch_reg,
        ins1_old_preg,
        ins1_new_preg,
        ins1_excp_code,
        ins1_excp_valid,
        ins1_special,
        ins1_is_store,
        ins1_valid
      },
      full,
      packet_pop,
      {
        cpacket_pc,
        cins0_register_allocated,
        cins0_arch_reg,
        cins0_old_preg,
        cins0_new_preg,
        cins0_excp_code,
        cins0_excp_valid,
        cins0_special,
        cins0_is_store,
        cins1_register_allocated,
        cins1_arch_reg,
        cins1_old_preg,
        cins1_new_preg,
        cins1_excp_code,
        cins1_excp_valid,
        cins1_special,
        cins1_is_store,
        cins1_valid
      },
      empty,
      rd_ptr,
      wr_ptr
  );
  assign rob0_status = {rd_ptr[3:0], 1'b0};
  assign rob1_status = {rd_ptr[3:0], 1'b1};
  assign rcu_pack = wr_ptr;
  //assign arch_reg0 = recoveryCounter0;
  //assign arch_reg1 = recoveryCounter1;
  assign sqb_commit0 = cins0_is_store & commit_ins0;
  assign sqb_commit1 = (cins1_is_store & commit_ins1);

  assign altcommit0 = altcommit & !partial_retire;
  assign altcommit1 = altcommit & partial_retire;
  srmt architectural_register_map (
      cpu_clock_i,
      p0_logical_reg_i,
      p0_phys_reg_o,
      p1_logical_reg_i,
      p1_phys_reg_o,
      p2_logical_reg_i,
      p2_phys_reg_o,
      p3_logical_reg_i,
      p3_phys_reg_o,
      p4_logical_reg_i,
      p4_phys_reg_o,
      p5_logical_reg_i,
      p5_phys_reg_o,
      cins0_arch_reg,
      cins0_new_preg,
      (commit_ins0 | altcommit0) & (cins0_register_allocated) & (cins0_arch_reg != 0),
      cins1_arch_reg,
      cins1_new_preg,
      (commit_ins1 | altcommit1) & (cins1_register_allocated) & (cins1_arch_reg != 0)
  );

  assign rcu_busy = full|!(retire_control_state==Normal||retire_control_state==TakeInterrupt||retire_control_state==ReclaimAndRecover);
  wire [29:0] currentPC = cpacket_pc[0] ? cpacket_pc : {cpacket_pc[29:1], partial_retire};
  wire [29:0] pcPlus4 = currentPC + 30'd1;  // used in special types CSRRW, SFENCE, FENCE.I
  // Conditions of committing
  assign packet_pop = ((partial_retire&(commit_ins1|altcommit1))|((commit_ins0|altcommit0)&((!cins1_valid)|(commit_ins1))))|(retire_control_state==ReclaimAndRecover);
  assign wr_data0 = retire_control_state == ReclaimAndRecover ? cins0_new_preg : cins0_old_preg;
  assign wr_data1 = retire_control_state == ReclaimAndRecover ? cins1_new_preg : cins1_old_preg;
  assign wr_en0 = retire_control_state==Normal ? (cins0_register_allocated)&(commit_ins0|altcommit0)&!(cins0_old_preg==0) : (retire_control_state==ReclaimAndRecover)
    &&cins0_register_allocated&&!empty&&!partial_retire;
  assign wr_en1 = retire_control_state==Normal ? (cins1_register_allocated)&(commit_ins1|altcommit1)&!(cins1_old_preg==0) : (retire_control_state==ReclaimAndRecover)
    &&cins1_register_allocated&&!empty;
  assign flush_o = retire_control_state == ReclaimAndRecover;
  assign commit_ins0 = (rob0_status_i)&&!empty&&!partial_retire&&!(cins0_excp_valid)&&!(|cins0_special) && (retire_control_state==Normal) && ((rob0_status!=exception_rob[4:0])||!exception_valid) && !rcu_block;
  assign commit_ins1 = (partial_retire|commit_ins0) && ((rob1_status_i)&&!empty&&!(cins1_excp_valid)&&!(|cins1_special)) && (retire_control_state==Normal) && ((rob1_status!=exception_rob[4:0])||!exception_valid) && !rcu_block && cins1_valid;
  wire older_alu = exception_rob[5]==rob_i[5] ? rob_i[4:0] < exception_rob[4:0] : rob_i[4:0] > exception_rob[4:0];
  wire oldest_live_excp = !exception_i ? 1'b0: !alu_excp_i ? 1'b1 : completed_rob_id[5]==rob_i[5] ? completed_rob_id[4:0]<rob_i[4:0] :
    completed_rob_id[4:0]>rob_i[4:0]; // 1 when LSU is oldest
  wire [5:0] winner = oldest_live_excp ? completed_rob_id : rob_i;
  wire older_than_current = (!exception_valid||(exception_rob[5]==winner[5] ? winner[4:0]<exception_rob[4:0] : winner[4:0]>exception_rob[4:0]))
    &&(alu_excp_i|exception_i); // 1 when older than current
  always_ff @(posedge cpu_clock_i) begin
    exception_valid <= rename_flush_o ? 1'b0 : exception_valid | (alu_excp_i | exception_i);
    exception_code <= older_than_current ? oldest_live_excp ? exception_code_i : alu_excp_code_i : exception_code;
    exception_rob <= older_than_current ? oldest_live_excp ? completed_rob_id : rob_i : exception_rob;
    relavant_address <= older_than_current & oldest_live_excp ? exception_addr : relavant_address;
    c1_btb_vpc <= (older_alu | !exception_valid) && alu_excp_i ? c1_btb_vpc_i : c1_btb_vpc;
    c1_btb_target <= (older_alu | !exception_valid) && alu_excp_i ? c1_btb_target_i : c1_btb_target;
    c1_cntr_pred <= (older_alu | !exception_valid) && alu_excp_i ? c1_cntr_pred_i : c1_cntr_pred;
    c1_bnch_tkn <= (older_alu | !exception_valid) && alu_excp_i ? c1_bnch_tkn_i : c1_bnch_tkn;
    c1_bnch_type <= (older_alu | !exception_valid) && alu_excp_i ? c1_bnch_type_i : c1_bnch_type;
    c1_bnch_present <=  (older_alu|!exception_valid)&&alu_excp_i ? c1_bnch_present_i : c1_bnch_present; /* Eliminate */
  end
  wire [3:0] int_type;
  wire       interrupt_pending;
  wire [3:0] excp_excp_code = partial_retire ? cins1_excp_code : cins0_excp_code;
  wire       excp_excp_valid = partial_retire ? cins1_excp_valid : cins0_excp_valid;
  wire [3:0] excp_special = partial_retire ? cins1_special : cins0_special;
  interrupt_router interrupts (
      cpm,
      mie,
      machine_interrupts,
      interrupt_pending,
      int_type
  );
  wire backendException = exception_valid && (partial_retire ? rob1_status==exception_rob[4:0] : rob0_status==exception_rob[4:0]) && !empty;
  reg altcommitted_on_interrupt = 0;
  reg [29:0] altcommit_npc = 0;
  assign oldest_instruction = {rd_ptr[3:0], partial_retire};
  assign rcu_block = retire_control_state != Normal && retire_control_state != ReclaimAndRecover;
  assign rename_flush_o = (retire_control_state==Await) && icache_idle && dcache_flush_resp && !mem_block_i;
  assign ins_commit0 = commit_ins0 | altcommit0;
  assign ins_commit1 = commit_ins1 | altcommit1;
  reg wfi = 0;
  assign mret = ((excp_special[2]))&(retire_control_state==Normal)&!empty&!mem_block_i&!excp_excp_valid;
  assign take_interrupt = retire_control_state == TakeInterrupt && !empty && !mem_block_i;
  assign take_exception = (excp_excp_valid|(backendException&!exception_code[4]))&!mem_block_i&!empty&(retire_control_state==Normal);
  assign tmu_epc_o = wfi ? pcPlus4 : altcommitted_on_interrupt ? altcommit_npc : currentPC;
  assign tmu_mcause_o = take_interrupt ? int_type : excp_excp_valid ? excp_excp_code : exception_code[3:0];
  assign tmu_mtval_o = backendException ? relavant_address : excp_excp_code[3:1]==0 ? {currentPC,2'b00} : 0;
  assign altcommit = ((backendException&exception_code[4])||((|excp_special)&&((excp_special[3]&(partial_retire ? rob1_status_i : rob0_status_i))||!excp_special[3])))
    && (retire_control_state==Normal)&!mem_block_i&!empty&!excp_special[0];
  reg btb_mod;

  // Special[3] == CSR writes
  // Special[2] == MRET (interrupts wont take place)
  // Special[1] == FENCE.I
  // Special[0] == WFI
  reg [3:0] retire_lim;
  always_ff @(posedge cpu_clock_i) begin
    case (retire_control_state)
      Normal: begin
        if (interrupt_pending&&(!empty)&&!mem_block_i&&((commit_ins0|commit_ins1|altcommit)|wfi)) begin
          retire_control_state <= TakeInterrupt;
          altcommit_npc <= (backendException & exception_code[4]) ? c1_btb_target : pcPlus4;
          altcommitted_on_interrupt <= altcommit;
          flush_address <= !(|mtvec_i[1:0]) ? mtvec_i[31:2] : {mtvec_i[31:2]} + {26'h0, tmu_mcause_o[3:0]};
        end else if ((excp_excp_valid | backendException) & !mem_block_i & !empty) begin
          retire_control_state <= Await;
          flush_address <= backendException & exception_code[4] ? c1_btb_target : mtvec_i[31:2];
        end else if ((((|excp_special)&&((excp_special[3]&(partial_retire ? rob1_status_i : rob0_status_i))||!excp_special[3])&!(wfi&excp_special[0]))&!mem_block_i&!empty)) begin
          retire_control_state <= excp_special[1] ? WipeInstructionCache : excp_special[0] ? WaitForInterrupt : Await;
          flush_address <= excp_special[2] ? mepc_i : pcPlus4;
        end
        partial_retire <= partial_retire ? partial_retire&!(commit_ins1|altcommit1) : ((commit_ins0)&!commit_ins1&cins1_valid)|(altcommit0&cins1_valid);
        btb_mod <= exception_code[4] & backendException;
      end
      WipeInstructionCache: begin
        if (icache_idle && sqb_empty) begin
          retire_control_state <= WipeDataCache;
        end
      end
      WaitForInterrupt: begin
        if (interrupt_pending && (!empty) && !mem_block_i) begin
          retire_control_state <= Normal;
          wfi <= 1;
        end
      end
      TakeInterrupt: begin
        if (!empty && !mem_block_i) begin
          retire_control_state <= Await;
          wfi <= 0;
        end
      end
      WipeDataCache: begin
        if (dcache_flush_resp && sqb_empty) begin
          retire_control_state <= Await;
        end
      end
      ReclaimAndRecover: begin
        wfi <= 0;
        partial_retire <= 0;
        altcommitted_on_interrupt <= 0;
        recoveryCounter0 <= recoveryCounter0 + 5'd2;
        recoveryCounter1 <= recoveryCounter1 + 5'd2;
        btb_mod <= 0;
        if ((rd_ptr[3:0] == retire_lim) || empty) begin
          retire_control_state <= Normal;
        end
      end
      Await: begin
        wfi <= 0;
        retire_lim <= wr_ptr[3:0] - 1'b1;
        if (icache_idle && dcache_flush_resp && !mem_block_i) begin
          retire_control_state <= ReclaimAndRecover;
        end
      end
      default: begin
        retire_control_state <= Normal;
      end
    endcase
  end
  assign icache_flush = icache_idle && sqb_empty && (retire_control_state == WipeInstructionCache);
  assign dcache_flush_o = dcache_flush_resp && sqb_empty && (retire_control_state == WipeDataCache);
  assign c1_btb_vpc_o = c1_btb_vpc;
  assign c1_btb_target_o = c1_btb_target;
  assign c1_cntr_pred_o = c1_cntr_pred;
  assign c1_bnch_tkn_o = c1_bnch_tkn;
  assign c1_bnch_type_o = c1_bnch_type;
  assign c1_btb_mod_o = (retire_control_state==Await)&&icache_idle&&dcache_flush_resp&&btb_mod&&!mem_block_i;
  assign c1_call_affirm_o = (rob0_call_i & commit_ins0) | (rob1_call_i & commit_ins1);
  assign c1_ret_affirm_o = (rob0_ret_i & commit_ins0) | (rob1_ret_i & commit_ins1);
endmodule
