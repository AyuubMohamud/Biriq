`define ALU_ADD 6'h00
`define ALU_SUB 6'h01
`define ALU_SLL 6'h02
`define ALU_SLT 6'h03
`define ALU_SLTU 6'h04
`define ALU_XOR 6'h08
`define ALU_SRL 6'h06
`define ALU_SRA 6'h07
`define ALU_OR 6'h09
`define ALU_AND 6'h0A
// Zba
`define ALU_SHXADD 6'h20
// Zbb
`define ALU_ANDN 6'h2A
`define ALU_ORN 6'h29
`define ALU_XNOR 6'h28
`define ALU_CTZ 6'h30
`define ALU_CLZ 6'h31
`define ALU_CPOP 6'h32
`define ALU_ROR 6'h26
`define ALU_ROL 6'h22
`define ALU_MAX 6'h34
`define ALU_MIN 6'h35
`define ALU_MAXU 6'h36
`define ALU_MINU 6'h37
`define ALU_SEXTB 6'h3C
`define ALU_SEXTH 6'h3D
`define ALU_ZEXTH 6'h3F
`define ALU_ORCB 6'h1B
`define ALU_REV8 6'h10
// Zbs
`define ALU_BEXT 6'h14
`define ALU_BCLR 6'h15
`define ALU_BINV 6'h16
`define ALU_BSET 6'h17
// Zbkb
`define ALU_PACK 6'h11
`define ALU_PACKH 6'h12
`define ALU_BREV8 6'h13
`define ALU_ZIP 6'h2C
`define ALU_UNZIP 6'h2D
// Zbkx
`define ALU_XPERM4 6'h2E
`define ALU_XPERM8 6'h2F
