module frontend #(
    parameter [31:0] C_START_ADDR = 32'h0,
    parameter [31:0] C_BPU_ENTRIES = 32,
    parameter C_BPU_ENABLE_RAS = 1,
    parameter C_BPU_RAS_ENTRIES = 32,
    parameter C_ICACHE_SIZE = 16384
) (
    input  wire logic        core_clock_i,
    input  wire logic        core_reset_i,
    input  wire logic        core_flush_i,
    input  wire logic [29:0] core_flush_pc,
    input  wire logic        enable_branch_pred,
    input  wire logic        enable_counter_overload,
    input  wire logic        counter_overload,
    input  wire logic        current_privlidge,
    input  wire logic        tw,
    input  wire logic [ 1:0] cbie,
    input  wire logic        cbcfe,
    input  wire logic        cbze,
    // System control port
    input  wire logic        cache_flush_i,
    // 00 - FLUSH, 01, Toggle ON/OFF, 1x undefined
    output wire logic        flush_resp_o,

    // TileLink Bus Master Uncached Heavyweight
    output logic      [ 2:0] icache_a_opcode,
    output logic      [ 2:0] icache_a_param,
    output logic      [ 3:0] icache_a_size,
    output logic      [31:0] icache_a_address,
    output logic      [ 3:0] icache_a_mask,
    output logic      [31:0] icache_a_data,
    output logic             icache_a_corrupt,
    output logic             icache_a_valid,
    input  wire logic        icache_a_ready,

    input  wire logic [ 2:0] icache_d_opcode,
    input  wire logic [ 1:0] icache_d_param,
    input  wire logic [ 3:0] icache_d_size,
    input  wire logic        icache_d_denied,
    input  wire logic [31:0] icache_d_data,
    input  wire logic        icache_d_corrupt,
    input  wire logic        icache_d_valid,
    output wire logic        icache_d_ready,
    // out to engine
    output logic             ins0_port_o,
    output logic             ins0_dnagn_o,
    output logic      [ 6:0] ins0_alu_type_o,
    output logic      [ 6:0] ins0_alu_opcode_o,
    output logic             ins0_alu_mc_o,
    output logic             ins0_alu_sc_o,
    output logic             ins0_alu_imm_o,
    output logic      [ 5:0] ins0_ios_type_o,
    output logic      [ 2:0] ins0_ios_opcode_o,
    output logic      [ 3:0] ins0_special_o,
    output logic      [ 4:0] ins0_rs1_o,
    output logic      [ 4:0] ins0_rs2_o,
    output logic      [ 4:0] ins0_dest_o,
    output logic      [31:0] ins0_imm_o,
    output logic      [ 2:0] ins0_reg_props_o,
    output logic             ins0_dnr_o,
    output logic             ins0_mov_elim_o,
    output logic      [ 1:0] ins0_hint_o,
    output logic             ins0_excp_valid_o,
    output logic      [ 3:0] ins0_excp_code_o,
    output logic             ins1_port_o,
    output logic             ins1_dnagn_o,
    output logic      [ 6:0] ins1_alu_type_o,
    output logic      [ 6:0] ins1_alu_opcode_o,
    output logic             ins1_alu_mc_o,
    output logic             ins1_alu_sc_o,
    output logic             ins1_alu_imm_o,
    output logic      [ 5:0] ins1_ios_type_o,
    output logic      [ 2:0] ins1_ios_opcode_o,
    output logic      [ 3:0] ins1_special_o,
    output logic      [ 4:0] ins1_rs1_o,
    output logic      [ 4:0] ins1_rs2_o,
    output logic      [ 4:0] ins1_dest_o,
    output logic      [31:0] ins1_imm_o,
    output logic      [ 2:0] ins1_reg_props_o,
    output logic             ins1_dnr_o,
    output logic             ins1_mov_elim_o,
    output logic      [ 1:0] ins1_hint_o,
    output logic             ins1_excp_valid_o,
    output logic      [ 3:0] ins1_excp_code_o,
    output logic             ins1_valid_o,
    output logic      [29:0] insbundle_pc_o,
    output logic      [ 1:0] btb_btype_o,
    output logic      [ 1:0] btb_bm_pred_o,
    output logic      [29:0] btb_target_o,
    output logic             btb_vld_o,
    output logic             btb_idx_o,
    output logic             btb_way_o,
    output logic             valid_o,
    input  wire logic        rn_busy_i,

    input wire logic [29:0] c1_btb_vpc_i,
    input wire logic [29:0] c1_btb_target_i,
    input wire logic [ 1:0] c1_cntr_pred_i,
    input wire logic        c1_bnch_tkn_i,
    input wire logic [ 1:0] c1_bnch_type_i,
    input wire logic        c1_btb_mod_i,
    input wire logic        c1_btb_way_i,
    input wire logic        c1_btb_bm_i,
    input wire logic        c1_call_affirm_i,
    input wire logic        c1_ret_affirm_i,

    output wire logic [29:0] i_addr,
    input  wire logic        i_kill
);

endmodule
