.C_RESET_ADDR(C_RESET_ADDR)
.C_BPU_ENTRIES(C_BPU_ENTRIES)
.C_BPU_ENABLE_RAS(C_BPU_ENABLE_RAS)
.C_BPU_RAS_ENTRIES(C_BPU_RAS_ENTRIES)
.C_HARTID(C_HARTID)
.C_SQ_ENTRIES(C_SQ_ENTRIES)
.C_PMP_ENTRIES(C_PMP_ENTRIES)
.C_ITIM_SIZE(C_ITIM_SIZE)
.C_ICACHE_SIZE(C_ICACHE_SIZE)
.C_DTIM_SIZE(C_DTIM_SIZE)
.C_DCACHE_SIZE(C_DCACHE_SIZE)
.C_HAS_IOASSIST(C_HAS_IOASSIST)
.C_ITLB_ENTRIES(C_ITLB_ENTRIES)
.C_DTLB_ENTRIES(C_DTLB_ENTRIES)
.C_HAS_SUPERVISOR(C_HAS_SUPERVISOR)
.C_HAS_USER(C_HAS_USER)
.C_HAS_ZMMUL(C_HAS_ZMMUL)
.C_HAS_DIV(C_HAS_DIV)
.C_HAS_ZAAMO(C_HAS_ZAAMO)
.C_HAS_ZALRSC(C_HAS_ZALRSC)
.C_HAS_ZBA(C_HAS_ZBA)
.C_HAS_ZBB(C_HAS_ZBB)
.C_HAS_ZBS(C_HAS_ZBS)
.C_HAS_ZBKB(C_HAS_ZBKB)
.C_HAS_ZBKX(C_HAS_ZBKX)
