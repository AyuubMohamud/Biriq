module ifu (
    
);
    
endmodule
