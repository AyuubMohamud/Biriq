parameter [31:0] C_RESET_ADDR = 32'h0,

parameter [31:0] C_BPU_ENTRIES = 64,

parameter C_BPU_ENABLE_RAS = 1,

parameter C_BPU_RAS_ENTRIES = 8,

parameter C_HARTID = 0,

parameter C_SQ_ENTRIES = 8,

parameter C_PMP_ENTRIES = 4,

parameter C_ITIM_SIZE = 0,

parameter C_ICACHE_SIZE = 0,

parameter C_DTIM_SIZE = 0,

parameter C_DCACHE_SIZE = 0,

parameter C_HAS_IOASSIST = 0,

parameter C_ITLB_ENTRIES = 0,

parameter C_DTLB_ENTRIES = 0,

parameter C_HAS_SUPERVISOR = 0,

parameter C_HAS_USER = 0,

parameter C_HAS_ZMMUL = 0,

parameter C_HAS_DIV = 0,

parameter C_HAS_ZAAMO = 0,

parameter C_HAS_ZALRSC = 0,

parameter C_HAS_ZBA = 1,

parameter C_HAS_ZBB = 1,

parameter C_HAS_ZBS = 1,

parameter C_HAS_ZBKB = 0,

parameter C_HAS_ZBKX = 0
