module mrq (
    
);
    
endmodule
